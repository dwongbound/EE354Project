`timescale 1ns / 1ps

module vga_controller(
	input clk, //this clock must be a slow enough clock to view the changing positions of the objects
	input bright,
	input rst,
	input up, down, left, right,
	input [9:0] hCount, vCount, // Is iterated through the screen pixel by pixel to show content
	output reg [11:0] rgb,
	input [15:0] v_counter,
	input [4:0] tilt_intensity, // this only goes from 1 to 8
	// these two values dictate the center of the doodle, incrementing and decrementing them leads the block to move in certain directions
	output [15:0] xpos, ypos,
	input q_Done, q_I, q_Up, q_Down,
	output [7:0] up_count,
	output [3:0] vert_speed, // how many pixels it moves up or down per clock
	input [9:0] JUMP_HEIGHT,
	input is_in_middle,
	output [15:0] true_y // the y location without scrolling effect
);

    // Temp size of doodle's radius
    localparam DOODLE_RADIUS = 13;
	localparam DOODLE_LENGTH = 27;
	localparam PLAT_RADIUS_W = 32; // Width radius of platform
	localparam PLAT_RADIUS_H = 7; // Height radius of platform
	reg last_direction = 1;
	reg down_flag = 0; // Used to reset up_count
    
	// Temp variable used to calculate location of filled block
	wire block_fill;

	// Temp vars
	reg [15:0] temp_x = 406, temp_y = 477;
	reg [7:0] temp_up_count = 0; // To count how many pixels it went up
	reg [3:0] temp_vert_speed = 0;
	reg [15:0] temp_true_y = 477;

	// Const color values
	parameter BLACK = 12'b0000_0000_0000;
	parameter OFF_WHITE = 12'hFFC;
	parameter RED   = 12'b1111_0000_0000;
	parameter PINK = 12'hFDF;

	// Sprite to register. Since VGA is 12 bit, 4 bits per rgb
	// Notice by indexing rules, it's right_down_img[y][x] gives you correct value
	reg [11:0] right_down_img[DOODLE_LENGTH][DOODLE_LENGTH] = '{
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hed5,12'hed5,12'h000,12'hed5,12'hed5,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
		'{12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hed5,12'h000},
		'{12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hed5,12'hed5,12'h000},
		'{12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hed5,12'h000},
		'{12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
		'{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h684,12'h684,12'h684,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'h000,12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'h000,12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc}};

	reg [11:0] left_down_img[DOODLE_LENGTH][DOODLE_LENGTH] = '{
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hed5,12'hed5,12'h000,12'hed5,12'hed5,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000},
		'{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000},
		'{12'h000,12'hed5,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000},
		'{12'h000,12'hed5,12'hed5,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000},
		'{12'h000,12'hed5,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000},
		'{12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'h000,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'hed5,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h684,12'h684,12'h684,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000,12'h000},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h684,12'h000,12'h000,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc}};
	
	reg [11:0] platform[15][65] = '{
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h443,12'h000,12'h000,12'h443,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'h443,12'h443,12'h000,12'had7,12'had7,12'hcea,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'h443,12'h443,12'had7,12'had7,12'hcea,12'hcea,12'hcea,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h000,12'h000,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'h443,12'had7,12'hcea,12'hcea,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h000},
		'{12'hffc,12'hffc,12'h443,12'had7,12'had7,12'h7b3,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h000},
		'{12'hffc,12'h443,12'hcea,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'had7,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'h000},
		'{12'hffc,12'h000,12'hcea,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'had7,12'had7,12'had7,12'h7b3,12'had7,12'h7b3,12'had7,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'h000},
		'{12'h000,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'had7,12'h7b3,12'had7,12'h7b3,12'had7,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'h7b3,12'had7,12'h7b3,12'had7,12'had7,12'had7,12'had7,12'had7,12'h7b3,12'h7b3,12'h000},
		'{12'h000,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'had7,12'had7,12'h7b3,12'had7,12'h7b3,12'had7,12'had7,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'had7,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'had7,12'h7b3,12'h7b3,12'h000,12'h000},
		'{12'h000,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'had7,12'h7b3,12'h7b3,12'h000,12'h000,12'hffc},
		'{12'h000,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'had7,12'h7b3,12'h7b3,12'h7b3,12'h000,12'h000,12'hffc},
		'{12'hffc,12'h000,12'h000,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h000,12'h000,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'h000,12'h000,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h7b3,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'h000,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc}};

	reg [11:0] game_over[150][315] = '{
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hffc,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hffc,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hffc,12'hffc,12'hffc,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'h112,12'h112,12'h112,12'h112,12'h112,12'h112,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00},
		'{12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00,12'hf00}};

	reg [11:0] title[150][250] = '{
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfee,12'hfee,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hdaa,12'hc44,12'hc44,12'hd88,12'hffe,12'hfee,12'hfed,12'hfee,12'hfee,12'hffe,12'hfed,12'ha00,12'ha00,12'ha00,12'hecb,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfed,12'hb33,12'ha00,12'ha00,12'hb22,12'hfee,12'hfee,12'hfed,12'hfee,12'hfee,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'hc66,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfed,12'hb11,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfed,12'hfee,12'hffe,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hfed,12'hfee,12'hffe,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'hb33,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfed,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'hdaa,12'hffe,12'hfed,12'hfee,12'hfee,12'hffe,12'hd88,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfed,12'hffe,12'hfee,12'hfee,12'hfed,12'hecc,12'hecb,12'hecb,12'hecb,12'hecb,12'hedd,12'hfed,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfed,12'hb33,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hfed,12'hfee,12'hffe,12'hffe,12'hfed,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfec,12'hfee,12'hebb,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hffe,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hfed,12'hfee,12'hffe,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'hb11,12'hedd,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hedd,12'hecb,12'hecc,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hedd,12'hc76,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'heba,12'hffe,12'hffe,12'hffe,12'hffe},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfed,12'hfee,12'hfed,12'hc55,12'ha00,12'ha00,12'ha00,12'hb11,12'hfed,12'hedc,12'hfed,12'hfed,12'hfed,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'hecb,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfed,12'hc66,12'ha00,12'ha00,12'ha00,12'hc44,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfed,12'hfed,12'hedc,12'hfed,12'hfee,12'hfee,12'hfee,12'hfed,12'hfed,12'hfee,12'hfee,12'hebb,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hecb,12'hfee,12'hfee,12'hfee},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfed,12'hfed,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'hecc,12'hfec,12'hfed,12'hfed,12'hfed,12'hfed,12'hb33,12'ha00,12'ha00,12'ha00,12'hebb,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedb,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedb,12'hdaa,12'hd88,12'hd88,12'hd88,12'hecc,12'hfed,12'hfed,12'hfdc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hecc,12'hfed,12'hfed},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'heba,12'hdaa,12'hdaa,12'hfed,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfed,12'hfee,12'hffe,12'hfee,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hfec,12'hfed,12'heba,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hecc,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hd77,12'hebb,12'hfee,12'hffe,12'hecb,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hfee},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hedc,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfed,12'heba,12'hd77,12'hd77,12'hd88,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfdc,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfee},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hedd,12'hdaa,12'heba,12'heba,12'hfee,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfdc,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hc76,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hedd,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfed,12'hfee,12'hffe,12'hffe,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hecb,12'hc76,12'hc66,12'hd77,12'hedd,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'hb11,12'hedd,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'heba,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hedd,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'heba,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hfed,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'hedd,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfee,12'hfee,12'hfec,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hffe,12'hfed,12'hecc,12'hd88,12'hd77,12'hd88,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffe,12'hffe,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hfed,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'hedd,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hffe,12'hb22,12'ha00,12'ha00,12'ha00,12'hc55,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hecb,12'hdaa,12'hecc,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hd77,12'ha00,12'ha00,12'ha00,12'hd88,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hedb,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hffe,12'hffe,12'hffe,12'hffe,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfed,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hc66,12'ha00,12'ha00,12'ha00,12'hecb,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hffe,12'hc55,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hffe,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'hc55,12'hedd,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hd77,12'ha00,12'ha00,12'ha00,12'hb33,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hedc,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hb33,12'ha00,12'ha00,12'ha00,12'hedd,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfed,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'hd77,12'hedb,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hffe,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'hfdc,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hedd,12'hecc,12'hecb,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfed,12'hdaa,12'ha00,12'ha00,12'ha00,12'hb11,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfec,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hb33,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'hc44,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hdaa,12'hb11,12'ha00,12'ha00,12'hc76,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfed,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hedc,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hfee,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfee,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfec,12'hfed,12'hd77,12'ha00,12'ha00,12'ha00,12'hb22,12'hedb,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfdc,12'hfec,12'hfec,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'hd88,12'hedc,12'hfdc,12'hfec,12'hfec,12'hedc,12'hc44,12'ha00,12'ha00,12'ha00,12'hc66,12'hfdc,12'hedb,12'hedc,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfec,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfec,12'hfed,12'hfdc,12'hfec,12'hfec,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hedc,12'hfdc,12'hfdc,12'hfec,12'hfec,12'hfec,12'hfec,12'hfec,12'hfec,12'hfdc,12'hedc,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hfec,12'hfec,12'hfec,12'hfec,12'hedc,12'hedb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfec,12'hfec,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfdc,12'hfdc,12'hfec,12'hfec,12'hfdc,12'hd77,12'ha00,12'ha00,12'ha00,12'hb33,12'hedc,12'hfec,12'hfec,12'hedc,12'hfec,12'hfdc,12'hc76,12'ha00,12'ha00,12'ha00,12'hc66,12'hedc,12'hfec,12'hedc,12'hedc,12'hfec,12'hfdc,12'hfec,12'hfec,12'hedc,12'hfec,12'hedc,12'hb33,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'hedb,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hfed,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hfed,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hffe,12'hfee,12'hffe,12'hfdc,12'hfee,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfee,12'hffe,12'hedd,12'hb11,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'hb33,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hd99,12'ha00,12'ha00,12'ha00,12'hb11,12'hfed,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hfed,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfec,12'hfee,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'hdaa,12'hffe,12'hffe,12'hffe,12'hfee,12'hedc,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hfee,12'hfee,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'hb33,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hc66,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hfed,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hfee,12'hecc,12'heba,12'hd99,12'hd77,12'hd77,12'hd77,12'hd77,12'hdaa,12'heba,12'hebb,12'hedd,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'hd88,12'hffe,12'hffe,12'hffe,12'hffe,12'hedc,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hd77,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hfed,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'ha00,12'ha00,12'ha00,12'hb11,12'hfee,12'hfec,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hd99,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hd99,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfed,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hd88,12'hffe,12'hffe,12'hfee,12'hfee,12'hfdc,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hd77,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'hfee,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hedd,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfee,12'hffe,12'hffe,12'hffe,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'hd88,12'hffe,12'hffe,12'hffe,12'hfee,12'hfdc,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hffe,12'hffe,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hd88,12'hebb,12'heba,12'hd88,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd88},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hedc,12'hedd,12'hedd,12'hedd,12'hedd,12'hfed,12'hffe,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'hfee,12'hfed,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hffe,12'hffe,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfed,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'hd88,12'hffe,12'hffe,12'hfee,12'hfee,12'hedc,12'hffe,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hb11,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hfed,12'hfed,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hecc,12'hc55,12'hb22,12'hb11,12'ha00,12'ha00,12'hb11,12'hb22,12'hc55,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'hfee,12'hfed,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hd88,12'hdaa,12'heba,12'hdaa,12'hc66,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hfee,12'hfee,12'hfee,12'hfec,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hfee,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hc66,12'hfee,12'hfee,12'hffe,12'hfee,12'hffe,12'hecc,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfed,12'hfee},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hc55,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hebb,12'hc55,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hc76,12'hebb,12'hfee,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedd,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'hd88,12'hfed,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hecb,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hffe,12'hb22,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hffe,12'hfee,12'hffe,12'hfec,12'hffe,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hffe,12'hffe,12'hffe,12'hb33,12'ha00,12'ha00,12'ha00,12'hc66,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'hb33,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hc55,12'hebb,12'hfee,12'hfee,12'hfee},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'hb11,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hedd,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'hc55,12'hfed,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hedc,12'hffe,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hffe,12'hffe,12'hffe,12'hb33,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hebb,12'hfed,12'hedd,12'hedd,12'hedd,12'hedd,12'hedd,12'hedc,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hd99,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hd77,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'hb11,12'hfed,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hedc,12'hfee,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hffe,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hecb,12'hc44,12'hb33,12'hb33,12'hebb,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'hd77,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfec,12'hedb,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedc,12'hedc,12'hedc,12'hedb,12'hecb,12'hebb,12'hebb,12'hebb,12'hebb,12'hecb,12'hedc,12'hedc,12'hfec,12'hfdc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfdc,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hedc,12'hfdc,12'hedc,12'hecb,12'hb22,12'hb11,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hedc,12'hedc,12'hfdc,12'hedc,12'hedc,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hedb,12'hedc,12'hedc,12'hedc,12'hedc,12'hfdc,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hedc,12'hedc,12'hedc,12'hedb,12'hedb,12'hedb,12'hecb,12'hdaa,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedc,12'hfdc,12'hedc,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfdc,12'hedc,12'hedc,12'hedc,12'hfdc,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hecc,12'hfdc,12'hedc,12'hfdc,12'hedc,12'heba,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedb,12'hedc,12'hfec,12'hb11,12'ha00,12'ha00,12'ha00,12'hc44,12'hfdc,12'hedc,12'hedc,12'hd88,12'hb11,12'ha00,12'hb11,12'hecb,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hfec,12'hfdc,12'hedc,12'hedc,12'hfec,12'hc66,12'ha00,12'ha00,12'ha00,12'hb33,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hfdc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfed,12'hecb,12'hb33,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hd88,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfdc,12'hfed,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hb33,12'hc66,12'hecb,12'hebb,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfec,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'hb11,12'hd77,12'hc76,12'hc44,12'hb33,12'hb22,12'hb22,12'hb22,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfee,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'heba,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hedd,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hc44,12'hc55,12'hc44,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfdc,12'hfee,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hfee,12'hfee,12'hfed,12'hedd,12'hedd,12'hfed,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfdc,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'hb11,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hebb,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hecb,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfec,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hd99,12'hffe,12'hffe,12'hfed,12'hfed,12'hffe,12'hffe,12'hebb,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hecc,12'hfed,12'hffe,12'hfee,12'hfee,12'hfee,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hffe,12'hfed,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hedc,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hedd,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hffe,12'hb33,12'ha00,12'ha00,12'ha00,12'hdaa,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hecc,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hedc,12'hfee,12'hffe,12'hfed,12'hc76,12'hc66,12'hc76,12'hedd,12'hfee,12'hffe,12'hfee,12'hfec,12'hfed,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'hb11,12'hfed,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfed,12'hb11,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfec,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hfee,12'hfee,12'hfee,12'hfed,12'hfed,12'hffe,12'hfee,12'hffe,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hfed,12'hffe,12'hffe,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hfdc,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hedd,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'hd99,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfed,12'hfed,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfec,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfdc,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedc,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hb11,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hedd,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hdaa,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hedc,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hfee,12'hfee,12'hfee,12'hfed,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hedd,12'hb11,12'ha00,12'ha00,12'ha00,12'hb33,12'hfed,12'hffe,12'hffe,12'hffe,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfdc,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hb11,12'hb11,12'hb11,12'hc44,12'hc44,12'hc66,12'hc66,12'hd77,12'hd99,12'hecb,12'hfdc,12'hfed,12'hffe,12'hffe,12'hecc,12'heba,12'hebb,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hfee,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfed,12'hfed,12'hfee,12'hecc,12'hd99,12'hc76,12'hc44,12'hb22,12'hb22,12'hb22,12'hb33,12'hc44,12'hc66,12'hdaa,12'hedd,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hfec,12'hb11,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hedd,12'heba,12'hc76,12'hc44,12'hb11,12'hb11,12'hc44,12'hd88,12'hecc,12'hc44,12'ha00,12'ha00,12'ha00,12'hb11,12'hfee,12'hffe,12'hffe,12'hffe,12'hffc,12'hffc,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hecb,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hedd,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hedc,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hecc,12'hffe,12'hffe,12'hfee,12'hfee,12'hfed,12'hfed,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hffe,12'hfee,12'hffe,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hffe,12'hffe,12'hfdc,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'hdaa,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hfdc,12'hfed,12'hedd,12'hc76,12'ha00,12'ha00,12'ha00,12'hd99,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfdc,12'hb33,12'ha00,12'ha00,12'ha00,12'heba,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hfee,12'hffe,12'hffe,12'hfee,12'hc76,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hecc,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfed,12'hfed,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hb11,12'ha00,12'ha00,12'ha00,12'hfed,12'hffe,12'hfee,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfdc,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hc55,12'ha00,12'ha00,12'ha00,12'hd99,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hfed,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfec,12'hd77,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfee,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfec,12'hc66,12'ha00,12'ha00,12'ha00,12'heba,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hfee,12'hffe,12'hfed,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfdc,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hffe,12'hffe,12'hfee,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hfed,12'hfed,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hfed,12'hffe,12'hfee,12'hfee,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hedc,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hc76,12'ha00,12'ha00,12'ha00,12'hd88,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hecb,12'hfee,12'hffe,12'hfee,12'hfee,12'hedd,12'heba,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hffe,12'hffe,12'hc76,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hfed,12'hd88,12'ha00,12'ha00,12'ha00,12'hd88,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffe,12'hffe,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hfee,12'hfee,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hfee,12'hfee,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'hedc,12'hffe,12'hfee,12'hfee,12'hecc,12'ha00,12'ha00,12'ha00,12'ha00,12'hecc,12'hfee,12'hedc,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'hd77,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hc55,12'hb22,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hfee,12'hffe,12'hd88,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hdaa,12'ha00,12'ha00,12'ha00,12'hc66,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hecc,12'hffe,12'hfed,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hffe,12'hffe,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfdc,12'hffe,12'hc76,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hffe,12'hfee,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'hb22,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfed,12'hfed,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hb22,12'ha00,12'ha00,12'ha00,12'hfdc,12'hfee,12'hfee,12'hfee,12'hfee,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hfdc,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfee,12'hffe,12'hffe,12'hffe,12'hecb,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hedd,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hd88,12'hedd,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hffe,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'hd77,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'heba,12'ha00,12'ha00,12'ha00,12'hc44,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hffe,12'hffe,12'hfee,12'hc44,12'ha00,12'ha00,12'ha00,12'hb11,12'hecc,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfdc,12'hfee,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hffe,12'hfee,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hffe,12'hfec,12'hfec,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hfdc,12'hffe,12'hffe,12'hffe,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfec,12'hffe,12'hfee,12'hfee,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfee,12'hffe,12'hfee,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'hb11,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hd88,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hd99,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hc76,12'ha00,12'ha00,12'ha00,12'hc76,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hecb,12'ha00,12'ha00,12'ha00,12'hc55,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hedb,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfed,12'hfed,12'hfed,12'hedc,12'hb22,12'ha00,12'ha00,12'ha00,12'hb22,12'hfdc,12'hfec,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfec,12'hfed,12'hfed,12'hfed,12'hedc,12'hfed,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hfed,12'hfec,12'hfed,12'hd88,12'ha00,12'ha00,12'ha00,12'hb33,12'hfed,12'hfed,12'hfed,12'hfec,12'hfed,12'hfed,12'hfdc,12'hedc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hc44,12'ha00,12'ha00,12'ha00,12'hb11,12'hedb,12'hfed,12'hfed,12'hfed,12'hfed,12'hedb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'heba,12'hfed,12'hfed,12'hfed,12'hd88,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd88,12'hfed,12'hfed,12'hfed,12'hfed,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfec,12'hfec,12'hfed,12'hecb,12'heba,12'hc76,12'hb22,12'hb11,12'hb11,12'hb11,12'hb22,12'hb33,12'hc76,12'heba,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hc66,12'ha00,12'ha00,12'ha00,12'hc76,12'hfed,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfec,12'hd99,12'hd77,12'hd88,12'hecb,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hfdc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfec,12'hfed,12'hfed,12'hfed,12'hc55,12'ha00,12'ha00,12'ha00,12'hc76,12'hfed,12'hfed,12'hfed,12'hedc,12'hb22,12'ha00,12'ha00,12'ha00,12'hc66,12'hfed,12'hfed,12'hfed,12'hfec,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hedc,12'hfed,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hfed,12'hfed,12'hfed,12'hfed,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfdc,12'hfed,12'hfed,12'hfed,12'hfed,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfdc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hd77,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hb11,12'ha00,12'ha00,12'ha00,12'hd88,12'hfed,12'hfed,12'hfed,12'hfed,12'hedc,12'hb22,12'ha00,12'ha00,12'ha00,12'hebb,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfdc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hfed,12'hc44,12'ha00,12'ha00,12'ha00,12'hd88,12'hfed,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hfee,12'hffe,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'hfee,12'hffe,12'hfee,12'hfee,12'hecb,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hfed,12'hfed,12'hfee,12'hfee,12'hfee,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hebb,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hedd,12'hb33,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hc76,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hb11,12'ha00,12'ha00,12'ha00,12'hedd,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hc66,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hfec,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hffe,12'hfee,12'hffe,12'hfed,12'hb22,12'ha00,12'ha00,12'ha00,12'hd77,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hfed,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffe,12'hffe,12'hfee,12'hedc,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hebb,12'hfee,12'hfee,12'hfee,12'hfed,12'hfed,12'hffe,12'hfee,12'hd99,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hfed,12'hfec,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hecb,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hebb,12'hfee,12'hecb,12'hc66,12'hc66,12'hc76,12'hfed,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'heba,12'hdaa,12'hebb,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hdaa,12'ha00,12'ha00,12'ha00,12'hb11,12'hfed,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hc66,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hfec,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hffe,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hdaa,12'hfee,12'hffe,12'hfed,12'hb33,12'ha00,12'ha00,12'ha00,12'hc44,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hd99,12'hffe,12'hffe,12'hffe,12'hffe,12'hfec,12'heba,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hd88,12'heba,12'heba,12'hd77,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfed,12'hfee,12'hfec,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hc55,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hc66,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hffe,12'hfee,12'hfee,12'hfed,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hc66,12'ha00,12'ha00,12'ha00,12'hb22,12'hfee,12'hfec,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hfee,12'hfee,12'hffe,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hdaa,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hfee,12'hfee,12'hffe,12'hfee,12'hffe,12'hfec,12'hfee,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hedd,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hedd,12'hebb,12'hecb,12'hecb,12'hecb,12'hecc,12'hedd,12'hffe,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfdc,12'hffe,12'hfee,12'hfee,12'hebb,12'hebb,12'hffe,12'hffe,12'hffe,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hedd,12'hfed,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hffe,12'hfed,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc44,12'hffe,12'hffe,12'hffe,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'heba,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'heba,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'hc76,12'hffe,12'hffe,12'hffe,12'hffe,12'hfee,12'hedc,12'hfee,12'hfee,12'heba,12'hc55,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hc76,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffe,12'hfed,12'hffe,12'hffe,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hfed,12'hb22,12'ha00,12'ha00,12'hb33,12'hd88,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfee,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'hd77,12'hfec,12'hfee,12'hfee,12'hfee,12'hffe,12'hffe,12'hffe,12'hc76,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hfed,12'hfee,12'hffe,12'hedd,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hc76,12'hebb,12'hfee,12'hfee,12'hfee,12'hecc,12'hc44,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hedc,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hedd,12'hc55,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'heba,12'hfee,12'hfee,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hecb,12'hffe,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hedd,12'hb11,12'ha00,12'ha00,12'ha00,12'hb11,12'hecb,12'hffe,12'hfee,12'hfee,12'hffe,12'hffe,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hfed,12'hffe,12'hffe,12'hffe,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hedd,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hedc,12'hfee,12'hffe,12'hfee,12'hffe,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hecc,12'hebb,12'hebb,12'hecb,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hd88,12'hfee,12'hfee,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hfee,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'hedd,12'hfee,12'hfee,12'hfee,12'hedd,12'hb22,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hedd,12'hffe,12'hffe,12'hffe,12'hfee,12'hd77,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc55,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfec,12'hfee,12'hffe,12'hffe,12'hfee,12'hffe,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hd99,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb11,12'hd88,12'hfee,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hfee,12'hebb,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb33,12'heba,12'hfee,12'hd99,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hb11,12'ha00,12'ha00,12'hb11,12'hedd,12'hffe,12'hffe,12'hffe,12'hfee,12'hffe,12'hedd,12'hd88,12'hb33,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hebb,12'hfed,12'hffe,12'hffe,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hdaa,12'hb33,12'ha00,12'ha00,12'ha00,12'hb11,12'hc76,12'hedd,12'hfec,12'hfee,12'hffe,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hfee,12'hfee,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hb22,12'hedd,12'hb22,12'ha00,12'ha00,12'hb11,12'hedd,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfed,12'hfed,12'hedd,12'heba,12'hd77,12'hc66,12'hc55,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfee,12'hfee,12'hfed,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfee,12'hfdc,12'hfed,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hedc,12'hedc,12'hecb,12'hb11,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hedb,12'hedb,12'hc55,12'ha00,12'ha00,12'hc44,12'hedc,12'hfdc,12'hedc,12'hedc,12'hedc,12'hedb,12'hedc,12'hedc,12'hedb,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedc,12'hedc,12'hedc,12'hedc,12'hedc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hfee,12'hffe,12'hffe,12'hedd,12'hc66,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'ha00,12'hc66,12'hedd,12'hfee,12'hfee,12'hecb,12'hedd,12'hedd,12'hfed,12'hffe,12'hffe,12'hffe,12'hfee,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hc66,12'hc44,12'hc44,12'hc44,12'hc44,12'hd88,12'hecc,12'hfee,12'hffe,12'hfee,12'hfee,12'hedb,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hedc,12'hfee,12'hfee,12'hffe,12'hffe,12'hfee,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hfdc,12'hfee,12'hfee,12'hffe,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc},
		'{12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc,12'hffc}};

	always@(posedge clk, posedge rst) 
	begin
		if (rst || q_I)
		begin 
			// rough values for above lowest block 
			temp_x <= 406;
			temp_y <= 477;
			temp_up_count <= 0; // default
			temp_vert_speed <= 0;
			down_flag <= 0;
			temp_true_y <= 477;
		end
		else if (clk) begin
			// Update acceleration
			if (temp_up_count <= 13) temp_vert_speed <= 4;
			else if (temp_up_count > 13 && temp_up_count <= 26) temp_vert_speed <= 4;
			else if (temp_up_count > 26 && temp_up_count <= 39) temp_vert_speed <= 3;
			else if (temp_up_count > 39 && temp_up_count <= 52) temp_vert_speed <= 3;
			else if (temp_up_count > 52 && temp_up_count <= 65) temp_vert_speed <= 3;
			else if (temp_up_count > 65 && temp_up_count <= 78) temp_vert_speed <= 2;
			else if (temp_up_count > 78 && temp_up_count <= 91) temp_vert_speed <= 2;
			else if (temp_up_count > 91 && temp_up_count <= 104) temp_vert_speed <= 2;
			else if (temp_up_count > 104 && temp_up_count <= 117) temp_vert_speed <= 1;
			else if (temp_up_count > 124) temp_vert_speed <= 1;

			/* Note that the top left of the screen does NOT correlate to vCount=0 and hCount=0. The display_controller.v file has the 
				synchronizing pulses for both the horizontal sync and the vertical sync begin at vcount=0 and hcount=0. Recall that after 
				the length of the pulse, there is also a short period called the back porch before the display area begins. So effectively, 
				the top left corner corresponds to (hcount,vcount)~(144,35). Which means with a 640x480 resolution, the bottom right corner 
				corresponds to ~(783,515).  
			*/
			if (right && !q_I) begin
				temp_x <= temp_x + tilt_intensity; //change the amount you increment to make the speed faster 
				last_direction <= 1;
				if(temp_x >= 775)
					temp_x <= 144;
			end
			else if (left && !q_I) begin
				temp_x <= temp_x - tilt_intensity;
				last_direction <= 0;
				if (temp_x <= 143)
					temp_x <= 774;
			end
			if (q_Up) begin // Second or for debugging
				// Doodle should only move if he is below the middle of the screen
				// If he's past the middle, everything else should move
				if (is_in_middle == 0)
					temp_y <= temp_y - vert_speed;
				temp_up_count <= temp_up_count + vert_speed;
				temp_true_y <= temp_true_y - vert_speed;
				if (down_flag) begin
					temp_up_count <= 0;
					down_flag <= 0;
				end
			end
			else if (q_Down) begin
				down_flag <= 1;
				temp_y <= temp_y + vert_speed;
				temp_true_y <= temp_true_y + vert_speed;
				temp_up_count <= temp_up_count - vert_speed;
				if (temp_up_count <= 4) // next clock should be at least -4.
					temp_up_count <= 0;
			end
		end
	end

	// Create Doodle's hitbox
	assign block_fill = vCount >= (temp_y-DOODLE_RADIUS) && vCount <= (temp_y+DOODLE_RADIUS) && hCount >= (temp_x-DOODLE_RADIUS) && hCount <= (temp_x+DOODLE_RADIUS); 
	
	always@ (*)
    	if (~bright)
			rgb = BLACK; // force black if not bright
		else if (rst)
			rgb = BLACK;
		// Game over
		else if (q_Done)
			// These values are calculated given starting offset
			if (hCount > 297 && hCount < 621 && vCount > 160 && vCount < 310)
				rgb = game_over[vCount-160][hCount-297];
			else
				rgb = RED;
		// Platforms
		else if (B1==1) // 288,208
			rgb = platform[vCount+PLAT_RADIUS_H-208-v_counter][hCount+PLAT_RADIUS_W-288];
		else if (B2==1) // 406,498
			rgb = platform[vCount+PLAT_RADIUS_H-498-v_counter][hCount+PLAT_RADIUS_W-406];
		else if (B3==1) // 632,338
			rgb = platform[vCount+PLAT_RADIUS_H-338-v_counter][hCount+PLAT_RADIUS_W-632];
		else if (B4==1) // 232,108
			rgb = platform[vCount+PLAT_RADIUS_H-108-v_counter][hCount+PLAT_RADIUS_W-232];
		else if (B5==1) // 288,478
			rgb = platform[vCount+PLAT_RADIUS_H-478-v_counter][hCount+PLAT_RADIUS_W-288];
		else if (B6==1) // 406,153
			rgb = platform[vCount+PLAT_RADIUS_H-153-v_counter][hCount+PLAT_RADIUS_W-406];
		else if (B8==1) // 232,338
			rgb = platform[vCount+PLAT_RADIUS_H-338-v_counter][hCount+PLAT_RADIUS_W-232];
		else if (B9==1) // 338,308
			rgb = platform[vCount+PLAT_RADIUS_H-308-v_counter][hCount+PLAT_RADIUS_W-338];
		else if (B10==1) // 432,368
			rgb = platform[vCount+PLAT_RADIUS_H-368-v_counter][hCount+PLAT_RADIUS_W-432];
		else if (B11==1) // 632, 80
			rgb = platform[vCount+PLAT_RADIUS_H-80-v_counter][hCount+PLAT_RADIUS_W-632];
		else if (B12==1) // 180, 20
			rgb = platform[vCount+PLAT_RADIUS_H-20-v_counter][hCount+PLAT_RADIUS_W-180];
		else if (B13==1) // 444, -100
			rgb = platform[vCount+PLAT_RADIUS_H-(-100)-v_counter][hCount+PLAT_RADIUS_W-444];
		// Doodle 
		else if (block_fill)
			if (last_direction == 1)
				rgb = right_down_img[vCount+DOODLE_RADIUS-ypos][hCount+DOODLE_RADIUS-xpos];
			else
				rgb = left_down_img[vCount+DOODLE_RADIUS-ypos][hCount+DOODLE_RADIUS-xpos];
		// title
		else if (q_I)
			if (hCount > 400 && hCount < 650 && vCount > 165 && vCount < 315)
				rgb = title[vCount-165][hCount-400];
			else
				rgb = OFF_WHITE;
		// Lines
		else if (vCount % 30 == 0)
			rgb = PINK;
		else
			rgb = OFF_WHITE; // background color

    assign B1 = (hCount >= (288-PLAT_RADIUS_W) && hCount <= (288+PLAT_RADIUS_W)) && (vCount>=(208-PLAT_RADIUS_H+v_counter) && vCount<=(208+PLAT_RADIUS_H+v_counter));
	assign B2 = (hCount >= (406-PLAT_RADIUS_W) && hCount <= (406+PLAT_RADIUS_W)) && (vCount>=(498-PLAT_RADIUS_H+v_counter) && vCount<=(498+PLAT_RADIUS_H+v_counter));
	assign B3 = (hCount >= (632-PLAT_RADIUS_W) && hCount <= (632+PLAT_RADIUS_W)) && (vCount>=(338-PLAT_RADIUS_H+v_counter) && vCount<=(338+PLAT_RADIUS_H+v_counter));
	assign B4 = (hCount >= (232-PLAT_RADIUS_W) && hCount <= (232+PLAT_RADIUS_W)) && (vCount>=(108-PLAT_RADIUS_H+v_counter) && vCount<=(108+PLAT_RADIUS_H+v_counter));
	assign B5 = (hCount >= (288-PLAT_RADIUS_W) && hCount <= (288+PLAT_RADIUS_W)) && (vCount>=(478-PLAT_RADIUS_H+v_counter) && vCount<=(478+PLAT_RADIUS_H+v_counter));
	assign B6 = (hCount >= (406-PLAT_RADIUS_W) && hCount <= (406+PLAT_RADIUS_W)) && (vCount>=(153-PLAT_RADIUS_H+v_counter) && vCount<=(153+PLAT_RADIUS_H+v_counter));
	assign B8 = (hCount >= (232-PLAT_RADIUS_W) && hCount <= (232+PLAT_RADIUS_W)) && (vCount>=(338-PLAT_RADIUS_H+v_counter) && vCount<=(338+PLAT_RADIUS_H+v_counter));
	assign B9 = (hCount >= (338-PLAT_RADIUS_W) && hCount <= (338+PLAT_RADIUS_W)) && (vCount>=(308-PLAT_RADIUS_H+v_counter) && vCount<=(308+PLAT_RADIUS_H+v_counter));
	assign B10 = (hCount >= (432-PLAT_RADIUS_W) && hCount <= (432+PLAT_RADIUS_W)) && (vCount>=(368-PLAT_RADIUS_H+v_counter) && vCount<=(368+PLAT_RADIUS_H+v_counter));
	assign B11 = (hCount >= (632-PLAT_RADIUS_W) && hCount <= (632+PLAT_RADIUS_W)) && (vCount>=(80-PLAT_RADIUS_H+v_counter) && vCount<=(80+PLAT_RADIUS_H+v_counter));
	assign B12 = (hCount >= (180-PLAT_RADIUS_W) && hCount <= (180+PLAT_RADIUS_W)) && (vCount>=(20-PLAT_RADIUS_H+v_counter) && vCount<=(20+PLAT_RADIUS_H+v_counter));
	assign B13 = (hCount >= (444-PLAT_RADIUS_W) && hCount <= (444+PLAT_RADIUS_W)) && (vCount>=((-100)-PLAT_RADIUS_H+v_counter) && vCount<=((-100)+PLAT_RADIUS_H+v_counter));
	
	// Assign temp vars to outputs
	assign xpos = temp_x;
	assign ypos = temp_y;
	assign up_count = temp_up_count;
	assign vert_speed = temp_vert_speed;
	assign true_y = temp_true_y;

endmodule